// 4 bits carry lookahead adder but returns c3 output.
module cla4_ov(a, b, ci, c3, co, s);
	input [3:0] a, b;
	input ci;
	output c3, co;
	output [3:0] s;
	
	wire c1, c2;
	
	fa_v2 u0_fa (.a(a[0]), .b(b[0]), .ci(ci), .s(s[0]));
	fa_v2 u1_fa (.a(a[1]), .b(b[1]), .ci(c1), .s(s[1]));
	fa_v2 u2_fa (.a(a[2]), .b(b[2]), .ci(c2), .s(s[2]));
	fa_v2 u3_fa (.a(a[3]), .b(b[3]), .ci(c3), .s(s[3]));
	clb4 u4_clb4 (.a(a), .b(b), .ci(ci), .c1(c1), .c2(c2), .c3(c3), .co(co));
endmodule
