module cla4(a, b, ci, co, s);
	input [3:0] a, b;
	input ci;
	output co;
	output [3:0] s;
	
	wire [2:0] c;
	
	fa_v2 u0_fa (.a(a[0]), .b(b[0]), .ci(ci), .s(s[0]));
	fa_v2 u1_fa (.a(a[1]), .b(b[1]), .ci(c[0]), .s(s[1]));
	fa_v2 u2_fa (.a(a[2]), .b(b[2]), .ci(c[1]), .s(s[2]));
	fa_v2 u3_fa (.a(a[3]), .b(b[3]), .ci(c[2]), .s(s[3]));
	clb4 u4_clb4 (.a(a), .b(b), .ci(ci), .c1(c[0]), .c2(c[1]), .c3(c[2]), .co(co));
	
endmodule
